// You can insert code here by setting file_header_inc in file execute_common.tpl

//=============================================================================
// Project  : generated_execute_tb
//
// File Name: execute_top_test_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Nov 12 21:15:16 2025
//=============================================================================
// Description: Test package for execute_top
//=============================================================================

`ifndef EXECUTE_TOP_TEST_PKG_SV
`define EXECUTE_TOP_TEST_PKG_SV

package execute_top_test_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import execute_in_pkg::*;
  import forward_pkg::*;
  import execute_out_pkg::*;
  import execute_top_pkg::*;

  `include "execute_top_test.sv"

endpackage : execute_top_test_pkg

`endif // EXECUTE_TOP_TEST_PKG_SV

