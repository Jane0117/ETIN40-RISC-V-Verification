// You can insert code here by setting file_header_inc in file execute_common.tpl

//=============================================================================
// Project  : generated_execute_tb
//
// File Name: execute_out_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Nov 12 21:15:16 2025
//=============================================================================
// Description: Package for agent execute_out
//=============================================================================

package execute_out_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;
  import common::*;


  `include "execute_out_execute_out_tx.sv"
  `include "execute_out_config.sv"
  `include "execute_out_driver.sv"
  `include "execute_out_monitor.sv"
  `include "execute_out_sequencer.sv"
  `include "execute_out_coverage.sv"
  `include "execute_out_agent.sv"
  `include "execute_out_seq_lib.sv"

endpackage : execute_out_pkg
