// You can insert code here by setting file_header_inc in file execute_common.tpl

//=============================================================================
// Project  : generated_execute_tb
//
// File Name: execute_in_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Nov 12 21:15:16 2025
//=============================================================================
// Description: Package for agent execute_in
//=============================================================================

package execute_in_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;


  `include "execute_in_execute_tx.sv"
  `include "execute_in_config.sv"
  `include "execute_in_driver.sv"
  `include "execute_in_monitor.sv"
  `include "execute_in_sequencer.sv"
  `include "execute_in_coverage.sv"
  `include "execute_in_agent.sv"
  `include "execute_in_seq_lib.sv"

endpackage : execute_in_pkg
