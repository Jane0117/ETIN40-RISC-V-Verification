// You can insert code here by setting file_header_inc in file .\common.tpl

//=============================================================================
// Project  : generated_alu_tb
//
// File Name: alu_top_test_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Oct 30 18:55:14 2025
//=============================================================================
// Description: Test package for alu_top
//=============================================================================

`ifndef ALU_TOP_TEST_PKG_SV
`define ALU_TOP_TEST_PKG_SV

package alu_top_test_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;
  import alu_top_pkg::*;

  `include "alu_top_test.sv"

endpackage : alu_top_test_pkg

`endif // ALU_TOP_TEST_PKG_SV

