// You can insert code here by setting file_header_inc in file .\common.tpl

//=============================================================================
// Project  : generated_alu_tb
//
// File Name: alu_top_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Oct 30 18:55:14 2025
//=============================================================================
// Description: Package for alu_top
//=============================================================================

package alu_top_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;

  `include "alu_top_config.sv"
  `include "alu_top_seq_lib.sv"
  `include "alu_top_env.sv"

endpackage : alu_top_pkg

