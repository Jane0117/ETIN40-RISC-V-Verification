`timescale 1ns / 1ps

import common::*;

module decode_execute_props;
    // Placeholder for FPV assertions. Bind or reference decode_execute_top here.
endmodule
